library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package YAY is
        type digit is array (0 to 5) of std_logic_vector(0 to 6);
end package;